`timescale 1ns / 1ps
//////////////////////////////////////////////////////////////////////////////////
// Company: 
// Engineer: 
// 
// Create Date: 2016/12/20 14:54:22
// Design Name: 
// Module Name: vga_controller
// Project Name: 
// Target Devices: 
// Tool Versions: 
// Description: 
// 
// Dependencies: 
// 
// Revision:
// Revision 0.01 - File Created
// Additional Comments:
// 
//////////////////////////////////////////////////////////////////////////////////

module Snake_Control(
         input wire clk_4Hz,
         input wire [1:0] mode,
         input wire up,
         input wire down,
         input wire right,
         input wire left,
         input wire [5:0] apple_x,
         input wire [5:0] apple_y,
         
         input wire [3:0] node, //��displayģ�鴫�������߽ڵ�λ��
         
         //output reg [35:0] zhuanwan,//��¼ת��Ǯ  �ߵĵڶ���λ��  ֻ��¼��ͷ�����жϷ���
         output reg [3:0] cubenum,//�÷֣����15 
         output wire [5:0] head_x,
         output wire [5:0] head_y,
         
         output reg [5:0] node_cube_x,
         output reg [5:0] node_cube_y
         
	 // output reg apple_status
    );
    reg [1:0] direct;//���������˶��ķ��� 
    reg [5:0] cube_x[15:0];
    reg [5:0] cube_y[15:0];
    
    assign head_x = cube_x[0];
    assign head_y = cube_y[0];
    
    parameter UP = 0;
    parameter DOWN = 1;
    parameter LEFT = 2;
    parameter RIGHT = 3;
//reg change_to_left,change_to_right,change_to_up,change_to_down;

    always @ ( node ) begin
        case(node)
            0: begin  node_cube_x = cube_x[0]; node_cube_y = cube_y[0]; end
            1: begin  node_cube_x = cube_x[1]; node_cube_y = cube_y[1]; end
            2: begin  node_cube_x = cube_x[2]; node_cube_y = cube_y[2]; end
            3: begin  node_cube_x = cube_x[3]; node_cube_y = cube_y[3]; end
            4: begin  node_cube_x = cube_x[4]; node_cube_y = cube_y[4]; end
            5: begin  node_cube_x = cube_x[5]; node_cube_y = cube_y[5]; end
            6: begin  node_cube_x = cube_x[6]; node_cube_y = cube_y[6]; end
            7: begin  node_cube_x = cube_x[7]; node_cube_y = cube_y[7]; end
            8: begin  node_cube_x = cube_x[8]; node_cube_y = cube_y[8]; end
            9: begin  node_cube_x = cube_x[9]; node_cube_y = cube_y[9]; end
            10: begin  node_cube_x = cube_x[10]; node_cube_y = cube_y[10]; end
            11: begin  node_cube_x = cube_x[11]; node_cube_y = cube_y[11]; end
            12: begin  node_cube_x = cube_x[12]; node_cube_y = cube_y[12]; end
            13: begin  node_cube_x = cube_x[13]; node_cube_y = cube_y[13]; end
            14: begin  node_cube_x = cube_x[14]; node_cube_y = cube_y[14]; end
            15: begin  node_cube_x = cube_x[15]; node_cube_y = cube_y[15]; end
            default : begin  node_cube_x = cube_x[0]; node_cube_y = cube_y[0]; end
        endcase
    end

   initial
        begin
            cube_x[0] <= 20;
            cube_y[0] <= 15;
            
            cube_x[1] <= 20;
            cube_y[1] <= 14;
            
            cube_x[2] <= 20;
            cube_y[2] <= 13;
        
            cube_x[3] <= 0;
            cube_y[3] <= 0;
            
            cube_x[4] <= 0;
            cube_y[4] <= 0;
            
            cube_x[5] <= 0;
            cube_y[5] <= 0;
            
            cube_x[6] <= 0;
            cube_y[6] <= 0;
            
            cube_x[7] <= 0;
            cube_y[7] <= 0;
            
            cube_x[8] <= 0;
            cube_y[8] <= 0;
            
            cube_x[9] <= 0;
            cube_y[9] <= 0;
            
            cube_x[10] <= 0;
            cube_y[10] <= 0;
            
            cube_x[11] <= 0;
            cube_y[11] <= 0;
            
            cube_x[12] <= 0;
            cube_y[12] <= 0;
            
            cube_x[13] <= 0;
            cube_y[13] <= 0;
            
            cube_x[14] <= 0;
            cube_y[14] <= 0;
            
            cube_x[15] <= 0;
            cube_y[15] <= 0;
        
            //zhuanwan <= 0;
            
            cubenum<=0;//�Ե�ƻ������
            direct<=DOWN;
           
        end

   wire button_plus;
   assign button_plus = ( up | down | left | right );

    always @ ( posedge button_plus ) //�޸���ͷ�˶�����
        begin
            if( up == 1 ) if( direct != UP && direct != DOWN)
                direct <= UP;
            if( down == 1)if( direct != UP && direct != DOWN)
                direct <= DOWN;
            if( left == 1) if( direct != LEFT && direct != RIGHT)
                direct <= LEFT;
            if( right == 1) if( direct != LEFT && direct != RIGHT)
                direct <= RIGHT;
            
            if(mode != 1) direct <= DOWN;    
            
        end

always@(posedge clk_4Hz)
    begin
          if( mode!=1 )
               begin
                cube_x[0] <= 20;
                cube_y[0] <= 15;
                
                cube_x[1] <= 20;
                cube_y[1] <= 14;
                
                cube_x[2] <= 20;
                cube_y[2] <= 13;
            
                cube_x[3] <= 0;
                cube_y[3] <= 0;
                
                cube_x[4] <= 0;
                cube_y[4] <= 0;
                
                cube_x[5] <= 0;
                cube_y[5] <= 0;
                
                cube_x[6] <= 0;
                cube_y[6] <= 0;
                
                cube_x[7] <= 0;
                cube_y[7] <= 0;
                
                cube_x[8] <= 0;
                cube_y[8] <= 0;
                
                cube_x[9] <= 0;
                cube_y[9] <= 0;
                
                cube_x[10] <= 0;
                cube_y[10] <= 0;
                
                cube_x[11] <= 0;
                cube_y[11] <= 0;
                
                cube_x[12] <= 0;
                cube_y[12] <= 0;
                
                cube_x[13] <= 0;
                cube_y[13] <= 0;
                
                cube_x[14] <= 0;
                cube_y[14] <= 0;
                
                cube_x[15] <= 0;
                cube_y[15] <= 0;
            
                //zhuanwan <= 0;
                
                cubenum<=0;//�Ե�ƻ������
               
          end
        if( mode==1 )
            begin
                  /**************************************************///�жϳ���
                  //ײǽ 
                  if((direct == UP && cube_y[0] == 1) | (direct==DOWN && cube_y[0] ==  28) | (direct==LEFT && cube_x[0] == 1) | (direct==RIGHT && cube_x[0] == 38))
                        cubenum<=15;
                   //ײ�Լ� 
                   else if((cube_y[0]==cube_y[1]&&cube_x[0]==cube_x[1])|
                            (cube_y[0]==cube_y[2]&&cube_x[0]==cube_x[2])|
                            (cube_y[0]==cube_y[3]&&cube_x[0]==cube_x[3]&&cubenum>0)|
                            (cube_y[0]==cube_y[4]&&cube_x[0]==cube_x[4]&&cubenum>1)|
                            (cube_y[0]==cube_y[5]&&cube_x[0]==cube_x[5]&&cubenum>2)|
                            (cube_y[0]==cube_y[6]&&cube_x[0]==cube_x[6]&&cubenum>3)|
                            (cube_y[0]==cube_y[7]&&cube_x[0]==cube_x[7]&&cubenum>4)|
                            (cube_y[0]==cube_y[8]&&cube_x[0]==cube_x[8]&&cubenum>5)|
                            (cube_y[0]==cube_y[9]&&cube_x[0]==cube_x[9]&&cubenum>6)|
                            (cube_y[0]==cube_y[10]&&cube_x[0]==cube_x[10]&&cubenum>7)|
                            (cube_y[0]==cube_y[11]&&cube_x[0]==cube_x[11]&&cubenum>8)|
                            (cube_y[0]==cube_y[12]&&cube_x[0]==cube_x[12]&&cubenum>9)|
                            (cube_y[0]==cube_y[13]&&cube_x[0]==cube_x[13]&&cubenum>10)|
                            (cube_y[0]==cube_y[14]&&cube_x[0]==cube_x[14]&&cubenum>11)|
                            (cube_y[0]==cube_y[15]&&cube_x[0]==cube_x[15]&&cubenum>12))
                                  cubenum<=15;
                   //���������
                   else 
                       begin
                       
                            cube_x[1]<=cube_x[0];
                            cube_y[1]<=cube_y[0];
                            
                            cube_x[2]<=cube_x[1];
                            cube_y[2]<=cube_y[1];
                            
                            cube_x[3]<=cube_x[2];
                            cube_y[3]<=cube_y[2];
                            
                            cube_x[4]<=cube_x[3];
                            cube_y[4]<=cube_y[3];
                            
                            cube_x[5]<=cube_x[4];
                            cube_y[5]<=cube_y[4];
                            
                            cube_x[6]<=cube_x[5];
                            cube_y[6]<=cube_y[5];
                            
                            cube_x[7]<=cube_x[6];
                            cube_y[7]<=cube_y[6];
                            
                            cube_x[8]<=cube_x[7];
                            cube_y[8]<=cube_y[7];
                            
                            cube_x[9]<=cube_x[8];
                            cube_y[9]<=cube_y[8];
                            
                            cube_x[10]<=cube_x[9];
                            cube_y[10]<=cube_y[9];
                            
                            cube_x[11]<=cube_x[10];
                            cube_y[11]<=cube_y[10];
                            
                            cube_x[12]<=cube_x[11];
                            cube_y[12]<=cube_y[11];
                            
                            cube_x[13]<=cube_x[12];
                            cube_y[13]<=cube_y[12];
                            
                            cube_x[14]<=cube_x[13];
                            cube_y[14]<=cube_y[13];
                            
                            cube_x[15]<=cube_x[14];
                            cube_y[15]<=cube_y[14];
                            
                            
                            case(direct)   //�ƶ���ͷ
                            UP:
                                 cube_y[0] <= cube_y[0] - 1;
                            DOWN:
                                 cube_y[0] <= cube_y[0] + 1;
                            LEFT:
                                 cube_x[0] <= cube_x[0] - 1;
                            RIGHT:
                                 cube_x[0] <= cube_x[0] + 1;
                            endcase
                            
                           
                            /**************************************************///�ж��Ƿ�Ե�ƻ��  
                            if(cube_x[0] == apple_x && cube_y[0] == apple_y)
                            begin
                                 cubenum <= cubenum + 1;
                            end
            
                       end 
            end
            
    end

endmodule
